module imm_gen (
    input  [31:0] instr,
    output reg [31:0] imm
);

    wire [6:0] opcode = instr[6:0];

    always @(*) begin
        case (opcode)
            // I-Type (ADDI, LW, JALR, etc.)
            7'b0010011, 7'b0000011, 7'b1100111, 7'b1110011: 
                imm = {{20{instr[31]}}, instr[31:20]};

            // S-Type (SW)
            7'b0100011: 
                imm = {{20{instr[31]}}, instr[31:25], instr[11:7]};

            // B-Type (BEQ, BNE)
            // Scrambled: imm[12], imm[10:5], imm[4:1], imm[11]
            7'b1100011: 
                imm = {{20{instr[31]}}, instr[7], instr[30:25], instr[11:8], 1'b0};

            // U-Type (LUI, AUIPC)
            // Just the top 20 bits, shifted up
            7'b0110111, 7'b0010111: 
                imm = {instr[31:12], 12'b0};

            // J-Type (JAL)
            // Scrambled: imm[20], imm[10:1], imm[11], imm[19:12]
            7'b1101111: 
                imm = {{12{instr[31]}}, instr[19:12], instr[20], instr[30:21], 1'b0};

            default: imm = 32'b0;
        endcase
    end

endmodule
